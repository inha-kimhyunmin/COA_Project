`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/11/18 22:24:41
// Design Name: 
// Module Name: reg_file
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module reg_file (
    input clk,
    input rst,

    // ?���??��?�� ?��?��?�� ?��?��
    input  [4:0] rs_idx,
    input  [4:0] rt_idx,
    input  [4:0] write_idx,  // mux?��?�� ?��?��?�� 목적�? ?��?��?��

    // ?���??��?�� ?���?
    input        RegWrite,
    input [31:0] write_data,

    // ?���??��?�� ?���?
    output [31:0] rs_data,
    output [31:0] rt_data
);

  // 32�? 32-bit ?���??��?��
  reg [31:0] regs[0:31];
  integer i;

  // 리셋 ?�� 모든 ?���??��?�� 0?���? 초기?��
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      for (i = 0; i < 32; i = i + 1)
        regs[i] <= 32'd0;
    end else if (RegWrite && write_idx != 0) begin
      regs[write_idx] <= write_data;
    end
  end

  // ?��기는 ?��?�� 조합 ?���? (read?�� 비동�?)
  assign rs_data = regs[rs_idx];
  assign rt_data = regs[rt_idx];

endmodule